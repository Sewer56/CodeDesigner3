.CDL    (      8   l      t   �   <          \  H   extern %thisaddr strToHex EE a0 EE a1 \s0 s1 s2     strLen  ���'  � �  �0 �-�� -�� -  2      -�@ #@       -   #�  !      � C0� B0 
 $#A  !    0 B$      7 B$
 $#a  !    0 c$      7 c$  "� #� & 1&��  �$  �{ �{  �{0 �{ �@ �'extern %thisaddr strLen EE a0   ���'  �-    ��
 `      �� `           �$ B$��       �{ � �'