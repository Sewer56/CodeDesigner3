.CDL    P      `   �      �   ,   �   �      �   $     (     0     L          d     extern %thisaddr test1 EE a0    test2   test3   test4   ���'  �                    �{ � �'extern %thisaddr test2  test3   test4   ���'  �              �{ � �'extern %thisaddr test3  test4   ���'  �        �{ � �'extern %thisaddr test4  ���'  �   4  �{ � �' 